module icache(addr,instr);
input [8:0] addr;
output [31:0] instr;

parameter MEM_SIZE = 512;
reg [31:0] memory [0:MEM_SIZE-1];

assign instr = memory[addr];

initial begin

memory[0]<=32'h20040000;
memory[1]<=32'h8c900000;
memory[2]<=32'h8c910004;
memory[3]<=32'h8c920008;
memory[4]<=32'h8c93000c;
memory[5]<=32'h8c940010;
memory[6]<=32'h8c950014;
memory[7]<=32'h8c960018;
memory[8]<=32'h8c97001c;
memory[9]<=32'h20050000;
memory[10]<=32'h3c068d00;
memory[11]<=32'h2007000a;
memory[12]<=32'h018dc026;
memory[13]<=32'h0309c026;
memory[14]<=32'h030ac026;
memory[15]<=32'h030bc026;
memory[16]<=32'h23190000;
memory[17]<=32'h201d0008;
memory[18]<=32'h001def00;
memory[19]<=32'h201c001b;
memory[20]<=32'h001ce600;
memory[21]<=32'h0290a026;
memory[22]<=32'h02b1a826;
memory[23]<=32'h02d2b026;
memory[24]<=32'h02f3b826;
memory[25]<=32'h10a700a8;
memory[26]<=32'h20a50001;
memory[27]<=32'h22990000;
memory[28]<=32'h0c000028;
memory[29]<=32'h23340000;
memory[30]<=32'h22b90000;
memory[31]<=32'h0c000028;
memory[32]<=32'h23350000;
memory[33]<=32'h22d90000;
memory[34]<=32'h0c000028;
memory[35]<=32'h23360000;
memory[36]<=32'h22f90000;
memory[37]<=32'h0c000028;
memory[38]<=32'h23370000;
memory[39]<=32'h0800003f;
memory[40]<=32'h00194582;
memory[41]<=32'h310803fc;
memory[42]<=32'h00194b82;
memory[43]<=32'h312903fc;
memory[44]<=32'h00195182;
memory[45]<=32'h314a03fc;
memory[46]<=32'h00195880;
memory[47]<=32'h316b03fc;
memory[48]<=32'h01044020;
memory[49]<=32'h01244820;
memory[50]<=32'h01445020;
memory[51]<=32'h01645820;
memory[52]<=32'h8d080200;
memory[53]<=32'h8d290200;
memory[54]<=32'h8d4a0200;
memory[55]<=32'h8d6b0200;
memory[56]<=32'h00084600;
memory[57]<=32'h00094c00;
memory[58]<=32'h000a5200;
memory[59]<=32'h0109c820;
memory[60]<=32'h032ac820;
memory[61]<=32'h032bc820;
memory[62]<=32'h03e00008;
memory[63]<=32'h200200ff;
memory[64]<=32'h00021400;
memory[65]<=32'h20430100;
memory[66]<=32'h00031a00;
memory[67]<=32'h2063ffff;
memory[68]<=32'h02824824;
memory[69]<=32'h0283a024;
memory[70]<=32'h02a25024;
memory[71]<=32'h02a3a824;
memory[72]<=32'h02c25824;
memory[73]<=32'h02c3b024;
memory[74]<=32'h02e26024;
memory[75]<=32'h02e3b824;
memory[76]<=32'h028aa026;
memory[77]<=32'h02aba826;
memory[78]<=32'h02ccb026;
memory[79]<=32'h02e9b826;
memory[80]<=32'h200200ff;
memory[81]<=32'h00021200;
memory[82]<=32'h204300ff;
memory[83]<=32'h00031c00;
memory[84]<=32'h206300ff;
memory[85]<=32'h02824824;
memory[86]<=32'h0283a024;
memory[87]<=32'h02a25024;
memory[88]<=32'h02a3a824;
memory[89]<=32'h02c25824;
memory[90]<=32'h02c3b024;
memory[91]<=32'h02e26024;
memory[92]<=32'h02e3b824;
memory[93]<=32'h028ba026;
memory[94]<=32'h02aca826;
memory[95]<=32'h02c9b026;
memory[96]<=32'h02eab826;
memory[97]<=32'h200200ff;
memory[98]<=32'h2003ffff;
memory[99]<=32'h00621822;
memory[100]<=32'h02824824;
memory[101]<=32'h0283a024;
memory[102]<=32'h02a25024;
memory[103]<=32'h02a3a824;
memory[104]<=32'h02c25824;
memory[105]<=32'h02c3b024;
memory[106]<=32'h02e26024;
memory[107]<=32'h02e3b824;
memory[108]<=32'h028ca026;
memory[109]<=32'h02a9a826;
memory[110]<=32'h02cab026;
memory[111]<=32'h02ebb826;
memory[112]<=32'h10a70041;
memory[113]<=32'h22990000;
memory[114]<=32'h0c00007e;
memory[115]<=32'h23340000;
memory[116]<=32'h22b90000;
memory[117]<=32'h0c00007e;
memory[118]<=32'h23350000;
memory[119]<=32'h22d90000;
memory[120]<=32'h0c00007e;
memory[121]<=32'h23360000;
memory[122]<=32'h22f90000;
memory[123]<=32'h0c00007e;
memory[124]<=32'h23370000;
memory[125]<=32'h080000b2;
memory[126]<=32'h200200ff;
memory[127]<=32'h00021c00;
memory[128]<=32'h00031200;
memory[129]<=32'h03224024;
memory[130]<=32'h03234824;
memory[131]<=32'h200200ff;
memory[132]<=32'h00021a00;
memory[133]<=32'h03235024;
memory[134]<=32'h332b00ff;
memory[135]<=32'h00094a00;
memory[136]<=32'h000a5400;
memory[137]<=32'h000b5e00;
memory[138]<=32'h00086040;
memory[139]<=32'h011dc024;
memory[140]<=32'h13000001;
memory[141]<=32'h019c6026;
memory[142]<=32'h00096840;
memory[143]<=32'h013dc024;
memory[144]<=32'h13000001;
memory[145]<=32'h01bc6826;
memory[146]<=32'h000a7040;
memory[147]<=32'h015dc024;
memory[148]<=32'h13000001;
memory[149]<=32'h01dc7026;
memory[150]<=32'h000b7840;
memory[151]<=32'h017dc024;
memory[152]<=32'h13000001;
memory[153]<=32'h01fc7826;
memory[154]<=32'h018dc026;
memory[155]<=32'h0309c026;
memory[156]<=32'h030ac026;
memory[157]<=32'h030bc026;
memory[158]<=32'h23190000;
memory[159]<=32'h01aec026;
memory[160]<=32'h030ac026;
memory[161]<=32'h030bc026;
memory[162]<=32'h0308c026;
memory[163]<=32'h0018c202;
memory[164]<=32'h0338c820;
memory[165]<=32'h01cfc026;
memory[166]<=32'h030bc026;
memory[167]<=32'h0308c026;
memory[168]<=32'h0309c026;
memory[169]<=32'h0018c402;
memory[170]<=32'h0338c820;
memory[171]<=32'h01ecc026;
memory[172]<=32'h0308c026;
memory[173]<=32'h0309c026;
memory[174]<=32'h030ac026;
memory[175]<=32'h0018c602;
memory[176]<=32'h0338c820;
memory[177]<=32'h03e00008;
memory[178]<=32'h00136e02;
memory[179]<=32'h00137200;
memory[180]<=32'h01cd6820;
memory[181]<=32'h21b90000;
memory[182]<=32'h0c000028;
memory[183]<=32'h232d0000;
memory[184]<=32'h00dd7024;
memory[185]<=32'h00063040;
memory[186]<=32'h11c00001;
memory[187]<=32'h00dc3026;
memory[188]<=32'h020d8026;
memory[189]<=32'h02068026;
memory[190]<=32'h02308826;
memory[191]<=32'h02519026;
memory[192]<=32'h02729826;
memory[193]<=32'h08000015;
memory[194]<=32'h080000c2;
memory[195]=32'h00000000;
memory[196]=32'h00000000;
memory[197]=32'h00000000;
memory[198]=32'h00000000;
memory[199]=32'h00000000;
memory[200]=32'h00000000;
memory[201]=32'h00000000;
memory[202]=32'h00000000;
memory[203]=32'h00000000;
memory[204]=32'h00000000;
memory[205]=32'h00000000;
memory[206]=32'h00000000;
memory[207]=32'h00000000;
memory[208]=32'h00000000;
memory[209]=32'h00000000;
memory[210]=32'h00000000;
memory[211]=32'h00000000;
memory[212]=32'h00000000;
memory[213]=32'h00000000;
memory[214]=32'h00000000;
memory[215]=32'h00000000;
memory[216]=32'h00000000;
memory[217]=32'h00000000;
memory[218]=32'h00000000;
memory[219]=32'h00000000;
memory[220]=32'h00000000;
memory[221]=32'h00000000;
memory[222]=32'h00000000;
memory[223]=32'h00000000;
memory[224]=32'h00000000;
memory[225]=32'h00000000;
memory[226]=32'h00000000;
memory[227]=32'h00000000;
memory[228]=32'h00000000;
memory[229]=32'h00000000;
memory[230]=32'h00000000;
memory[231]=32'h00000000;
memory[232]=32'h00000000;
memory[233]=32'h00000000;
memory[234]=32'h00000000;
memory[235]=32'h00000000;
memory[236]=32'h00000000;
memory[237]=32'h00000000;
memory[238]=32'h00000000;
memory[239]=32'h00000000;
memory[240]=32'h00000000;
memory[241]=32'h00000000;
memory[242]=32'h00000000;
memory[243]=32'h00000000;
memory[244]=32'h00000000;
memory[245]=32'h00000000;
memory[246]=32'h00000000;
memory[247]=32'h00000000;
memory[248]=32'h00000000;
memory[249]=32'h00000000;
memory[250]=32'h00000000;
memory[251]=32'h00000000;
memory[252]=32'h00000000;
memory[253]=32'h00000000;
memory[254]=32'h00000000;
memory[255]=32'h00000000;
memory[256]=32'h00000000;
memory[257]=32'h00000000;
memory[258]=32'h00000000;
memory[259]=32'h00000000;
memory[260]=32'h00000000;
memory[261]=32'h00000000;
memory[262]=32'h00000000;
memory[263]=32'h00000000;
memory[264]=32'h00000000;
memory[265]=32'h00000000;
memory[266]=32'h00000000;
memory[267]=32'h00000000;
memory[268]=32'h00000000;
memory[269]=32'h00000000;
memory[270]=32'h00000000;
memory[271]=32'h00000000;
memory[272]=32'h00000000;
memory[273]=32'h00000000;
memory[274]=32'h00000000;
memory[275]=32'h00000000;
memory[276]=32'h00000000;
memory[277]=32'h00000000;
memory[278]=32'h00000000;
memory[279]=32'h00000000;
memory[280]=32'h00000000;
memory[281]=32'h00000000;
memory[282]=32'h00000000;
memory[283]=32'h00000000;
memory[284]=32'h00000000;
memory[285]=32'h00000000;
memory[286]=32'h00000000;
memory[287]=32'h00000000;
memory[288]=32'h00000000;
memory[289]=32'h00000000;
memory[290]=32'h00000000;
memory[291]=32'h00000000;
memory[292]=32'h00000000;
memory[293]=32'h00000000;
memory[294]=32'h00000000;
memory[295]=32'h00000000;
memory[296]=32'h00000000;
memory[297]=32'h00000000;
memory[298]=32'h00000000;
memory[299]=32'h00000000;
memory[300]=32'h00000000;
memory[301]=32'h00000000;
memory[302]=32'h00000000;
memory[303]=32'h00000000;
memory[304]=32'h00000000;
memory[305]=32'h00000000;
memory[306]=32'h00000000;
memory[307]=32'h00000000;
memory[308]=32'h00000000;
memory[309]=32'h00000000;
memory[310]=32'h00000000;
memory[311]=32'h00000000;
memory[312]=32'h00000000;
memory[313]=32'h00000000;
memory[314]=32'h00000000;
memory[315]=32'h00000000;
memory[316]=32'h00000000;
memory[317]=32'h00000000;
memory[318]=32'h00000000;
memory[319]=32'h00000000;
memory[320]=32'h00000000;
memory[321]=32'h00000000;
memory[322]=32'h00000000;
memory[323]=32'h00000000;
memory[324]=32'h00000000;
memory[325]=32'h00000000;
memory[326]=32'h00000000;
memory[327]=32'h00000000;
memory[328]=32'h00000000;
memory[329]=32'h00000000;
memory[330]=32'h00000000;
memory[331]=32'h00000000;
memory[332]=32'h00000000;
memory[333]=32'h00000000;
memory[334]=32'h00000000;
memory[335]=32'h00000000;
memory[336]=32'h00000000;
memory[337]=32'h00000000;
memory[338]=32'h00000000;
memory[339]=32'h00000000;
memory[340]=32'h00000000;
memory[341]=32'h00000000;
memory[342]=32'h00000000;
memory[343]=32'h00000000;
memory[344]=32'h00000000;
memory[345]=32'h00000000;
memory[346]=32'h00000000;
memory[347]=32'h00000000;
memory[348]=32'h00000000;
memory[349]=32'h00000000;
memory[350]=32'h00000000;
memory[351]=32'h00000000;
memory[352]=32'h00000000;
memory[353]=32'h00000000;
memory[354]=32'h00000000;
memory[355]=32'h00000000;
memory[356]=32'h00000000;
memory[357]=32'h00000000;
memory[358]=32'h00000000;
memory[359]=32'h00000000;
memory[360]=32'h00000000;
memory[361]=32'h00000000;
memory[362]=32'h00000000;
memory[363]=32'h00000000;
memory[364]=32'h00000000;
memory[365]=32'h00000000;
memory[366]=32'h00000000;
memory[367]=32'h00000000;
memory[368]=32'h00000000;
memory[369]=32'h00000000;
memory[370]=32'h00000000;
memory[371]=32'h00000000;
memory[372]=32'h00000000;
memory[373]=32'h00000000;
memory[374]=32'h00000000;
memory[375]=32'h00000000;
memory[376]=32'h00000000;
memory[377]=32'h00000000;
memory[378]=32'h00000000;
memory[379]=32'h00000000;
memory[380]=32'h00000000;
memory[381]=32'h00000000;
memory[382]=32'h00000000;
memory[383]=32'h00000000;
memory[384]=32'h00000000;
memory[385]=32'h00000000;
memory[386]=32'h00000000;
memory[387]=32'h00000000;
memory[388]=32'h00000000;
memory[389]=32'h00000000;
memory[390]=32'h00000000;
memory[391]=32'h00000000;
memory[392]=32'h00000000;
memory[393]=32'h00000000;
memory[394]=32'h00000000;
memory[395]=32'h00000000;
memory[396]=32'h00000000;
memory[397]=32'h00000000;
memory[398]=32'h00000000;
memory[399]=32'h00000000;
memory[400]=32'h00000000;
memory[401]=32'h00000000;
memory[402]=32'h00000000;
memory[403]=32'h00000000;
memory[404]=32'h00000000;
memory[405]=32'h00000000;
memory[406]=32'h00000000;
memory[407]=32'h00000000;
memory[408]=32'h00000000;
memory[409]=32'h00000000;
memory[410]=32'h00000000;
memory[411]=32'h00000000;
memory[412]=32'h00000000;
memory[413]=32'h00000000;
memory[414]=32'h00000000;
memory[415]=32'h00000000;
memory[416]=32'h00000000;
memory[417]=32'h00000000;
memory[418]=32'h00000000;
memory[419]=32'h00000000;
memory[420]=32'h00000000;
memory[421]=32'h00000000;
memory[422]=32'h00000000;
memory[423]=32'h00000000;
memory[424]=32'h00000000;
memory[425]=32'h00000000;
memory[426]=32'h00000000;
memory[427]=32'h00000000;
memory[428]=32'h00000000;
memory[429]=32'h00000000;
memory[430]=32'h00000000;
memory[431]=32'h00000000;
memory[432]=32'h00000000;
memory[433]=32'h00000000;
memory[434]=32'h00000000;
memory[435]=32'h00000000;
memory[436]=32'h00000000;
memory[437]=32'h00000000;
memory[438]=32'h00000000;
memory[439]=32'h00000000;
memory[440]=32'h00000000;
memory[441]=32'h00000000;
memory[442]=32'h00000000;
memory[443]=32'h00000000;
memory[444]=32'h00000000;
memory[445]=32'h00000000;
memory[446]=32'h00000000;
memory[447]=32'h00000000;
memory[448]=32'h00000000;
memory[449]=32'h00000000;
memory[450]=32'h00000000;
memory[451]=32'h00000000;
memory[452]=32'h00000000;
memory[453]=32'h00000000;
memory[454]=32'h00000000;
memory[455]=32'h00000000;
memory[456]=32'h00000000;
memory[457]=32'h00000000;
memory[458]=32'h00000000;
memory[459]=32'h00000000;
memory[460]=32'h00000000;
memory[461]=32'h00000000;
memory[462]=32'h00000000;
memory[463]=32'h00000000;
memory[464]=32'h00000000;
memory[465]=32'h00000000;
memory[466]=32'h00000000;
memory[467]=32'h00000000;
memory[468]=32'h00000000;
memory[469]=32'h00000000;
memory[470]=32'h00000000;
memory[471]=32'h00000000;
memory[472]=32'h00000000;
memory[473]=32'h00000000;
memory[474]=32'h00000000;
memory[475]=32'h00000000;
memory[476]=32'h00000000;
memory[477]=32'h00000000;
memory[478]=32'h00000000;
memory[479]=32'h00000000;
memory[480]=32'h00000000;
memory[481]=32'h00000000;
memory[482]=32'h00000000;
memory[483]=32'h00000000;
memory[484]=32'h00000000;
memory[485]=32'h00000000;
memory[486]=32'h00000000;
memory[487]=32'h00000000;
memory[488]=32'h00000000;
memory[489]=32'h00000000;
memory[490]=32'h00000000;
memory[491]=32'h00000000;
memory[492]=32'h00000000;
memory[493]=32'h00000000;
memory[494]=32'h00000000;
memory[495]=32'h00000000;
memory[496]=32'h00000000;
memory[497]=32'h00000000;
memory[498]=32'h00000000;
memory[499]=32'h00000000;
memory[500]=32'h00000000;
memory[501]=32'h00000000;
memory[502]=32'h00000000;
memory[503]=32'h00000000;
memory[504]=32'h00000000;
memory[505]=32'h00000000;
memory[506]=32'h00000000;
memory[507]=32'h00000000;
memory[508]=32'h00000000;
memory[509]=32'h00000000;
memory[510]=32'h00000000;
memory[511]=32'h00000000;


end

endmodule
